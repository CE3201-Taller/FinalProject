module seven_decoder
(
);
endmodule