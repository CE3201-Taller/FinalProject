/* 
 *
 *
 * @file  controller.sv
 * @autor Luis Arturo Mora Granados
 * @date  14/10/2018
 */

module controller
(
     input logic         clk_i, rst_i,
     input logic [31:12] instr_i,
     input logic [3:0]   alu_flags_i,
    output logic [1:0]   reg_src_o,
    output logic         reg_write_o,
    output logic [1:0]   imm_src_o,
    output logic         alu_src_o,
    output logic [1:0]   alu_control_o
    output logic         mem_write_o, mem_to_reg_o, 
    output logic         pc_src_o
);

    logic [1:0] flag_write;
    logic       pc_src, reg_write, men_write;

    decoder dec(instr_i[27:26], instr_i[25:20], instr_i[15:12],
                flag_write, pc_src, reg_write, men_write,
                mem_to_reg_o, alu_src_o, imm_src_o, reg_src_o, alu_control_o);

    condlogic c(clk_i, rst_i, instr_i[31:28], alu_flags_i,
                flag_write, pc_src, reg_write, men_write,
                pc_src_o, reg_write_o, mem_write_o);
endmodule
