module display_decoder
(
	 input logic [31:0] data_i,
	output logic [6:0]  display_1_o, display_2_o, display_3_o
);
endmodule